//FU
/*

inputs:

output:
     
*/
module FU (wr_add);



endmodule